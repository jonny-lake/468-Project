module move_register(r1,r2);
input [31:0]r2;
output [31:0]r1;

assign r1 = r2;

endmodule