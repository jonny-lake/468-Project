module Add(A, B, Sum);
	input [3:0] A, B;
	output [4:0] Sum;

	assign Sum = A+B;
endmodule
