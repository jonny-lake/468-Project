module move_IMM(r1,n);
input [15:0]n;
output [31:0]r1;

assign r1 = n;

endmodule
